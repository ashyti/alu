library ieee;
use ieee.std_logic_1164.all;

package globals is
	type aluop is (
		ADDS,
		MULTI
	);
end globals;
